module architecture(input clk);
wire [63:0] d,e,Writedata,immediateout, RD1,RD2, Mux1output, ALUOut, DataOutput, shiftoutput,Mux10output;
wire [31:0] RD, PC, PCPlus4;
wire [31:0] branchaddress,PCinput;
wire [3:0] Control; 
wire [1:0] Aluop,MemtoReg;
wire [31:0]PCaddress;
//wire b;
MUX #(32)M9(PCaddress,ALUOut[31:0],jump,PCinput);
PCCounter P1(clk,PCinput,PC);
adder A1(PC,PCPlus4);
instructionmemory I1(PC,RD);
mainController M1(RD[6:0],ALUSrc, MemtoReg, RegWrite, MemRead, MemWrite, Branch,jump,Asel,Aluop);
Registerfile R1(clk,RegWrite,RD[19:15],RD[24:20],RD[11:7],Writedata,RD1,RD2);
immediategeneration S1(RD[31:0],immediateout);
MUX #(64)M4(RD2,immediateout,ALUSrc,Mux1output);
//MUX #(1)M9(1'bx,RD[30],RD[5],b);
ALUControl A3(Aluop,RD[30],RD[14:12],Control);
MUX #(64)M10(RD1,PC,Asel,Mux10output);
assign d = {{32{Mux10output[31]}},Mux10output[31:0]};
ALU A2(Control,d,Mux1output,ALUOut,Zero);
DataMemory D1(clk,MemWrite,MemRead,ALUOut,RD2,DataOutput);
assign e = {{32{PCPlus4[31]}},PCPlus4[31:0]};
MUX1 #(64)M2(ALUOut,DataOutput,e,MemtoReg,Writedata);
and Q1(andoutput,Branch,Zero);
shift S12(immediateout,shiftoutput);
add A23(PC,shiftoutput[31:0],branchaddress);
MUX #(32)M3(PCPlus4,branchaddress,andoutput,PCaddress);
endmodule
